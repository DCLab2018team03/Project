`ifndef _PITCH_DEFINE_SV_
`define _PITCH_DEFINE_SV_
// window size for time-stretching and pitch-shifting, if you change the window size,
// remember to modify the hanning coefficients below
parameter [9:0] WindowSize = 10'd1024;
parameter [8:0] H_s = 9'd512;
parameter [8:0] tolerance = 9'd512;
parameter [11:0] AnalysisFrameSize = 12'd2560;
// hanning window parameter 0~511 (to use 512~1023, just call the symetric part)
// format: unsigned, the first bit is preserverd (in case they are used to be signed),
//         the remaining represents the floating point of the coefficients
//         (no precise 1 occurs, so it's OK not to store the int part)
parameter signed [19:0] HANN_C [WindowSize-1:0] = {
20'b00000000000000000000,
20'b00000000000000000100,
20'b00000000000000010011,
20'b00000000000000101100,
20'b00000000000001001111,
20'b00000000000001111011,
20'b00000000000010110001,
20'b00000000000011110010,
20'b00000000000100111100,
20'b00000000000110010000,
20'b00000000000111101110,
20'b00000000001001010110,
20'b00000000001011000111,
20'b00000000001101000011,
20'b00000000001111001000,
20'b00000000010001010111,
20'b00000000010011110000,
20'b00000000010110010011,
20'b00000000011001000000,
20'b00000000011011110110,
20'b00000000011110110111,
20'b00000000100010000001,
20'b00000000100101010101,
20'b00000000101000110011,
20'b00000000101100011010,
20'b00000000110000001100,
20'b00000000110100000111,
20'b00000000111000001100,
20'b00000000111100011010,
20'b00000001000000110011,
20'b00000001000101010101,
20'b00000001001010000001,
20'b00000001001110110110,
20'b00000001010011110110,
20'b00000001011000111111,
20'b00000001011110010001,
20'b00000001100011101101,
20'b00000001101001010011,
20'b00000001101111000011,
20'b00000001110100111100,
20'b00000001111010111111,
20'b00000010000001001011,
20'b00000010000111100001,
20'b00000010001110000001,
20'b00000010010100101010,
20'b00000010011011011100,
20'b00000010100010011001,
20'b00000010101001011110,
20'b00000010110000101101,
20'b00000010111000000110,
20'b00000010111111101000,
20'b00000011000111010011,
20'b00000011001111001000,
20'b00000011010111000110,
20'b00000011011111001110,
20'b00000011100111011111,
20'b00000011101111111001,
20'b00000011111000011101,
20'b00000100000001001001,
20'b00000100001010000000,
20'b00000100010010111111,
20'b00000100011100001000,
20'b00000100100101011001,
20'b00000100101110110100,
20'b00000100111000011001,
20'b00000101000010000110,
20'b00000101001011111100,
20'b00000101010101111100,
20'b00000101100000000100,
20'b00000101101010010110,
20'b00000101110100110000,
20'b00000101111111010100,
20'b00000110001010000001,
20'b00000110010100110110,
20'b00000110011111110100,
20'b00000110101010111100,
20'b00000110110110001100,
20'b00000111000001100101,
20'b00000111001101000111,
20'b00000111011000110001,
20'b00000111100100100100,
20'b00000111110000100000,
20'b00000111111100100101,
20'b00001000001000110011,
20'b00001000010101001001,
20'b00001000100001100111,
20'b00001000101110001110,
20'b00001000111010111110,
20'b00001001000111110110,
20'b00001001010100110111,
20'b00001001100010000000,
20'b00001001101111010010,
20'b00001001111100101100,
20'b00001010001010001110,
20'b00001010010111111001,
20'b00001010100101101011,
20'b00001010110011100111,
20'b00001011000001101010,
20'b00001011001111110110,
20'b00001011011110001001,
20'b00001011101100100101,
20'b00001011111011001001,
20'b00001100001001110101,
20'b00001100011000101001,
20'b00001100100111100101,
20'b00001100110110101001,
20'b00001101000101110101,
20'b00001101010101001000,
20'b00001101100100100100,
20'b00001101110100000111,
20'b00001110000011110010,
20'b00001110010011100101,
20'b00001110100011011111,
20'b00001110110011100001,
20'b00001111000011101011,
20'b00001111010011111100,
20'b00001111100100010101,
20'b00001111110100110101,
20'b00010000000101011101,
20'b00010000010110001100,
20'b00010000100111000010,
20'b00010000111000000000,
20'b00010001001001000101,
20'b00010001011010010001,
20'b00010001101011100101,
20'b00010001111101000000,
20'b00010010001110100001,
20'b00010010100000001010,
20'b00010010110001111010,
20'b00010011000011110001,
20'b00010011010101101111,
20'b00010011100111110011,
20'b00010011111001111111,
20'b00010100001100010001,
20'b00010100011110101010,
20'b00010100110001001010,
20'b00010101000011110001,
20'b00010101010110011110,
20'b00010101101001010010,
20'b00010101111100001100,
20'b00010110001111001101,
20'b00010110100010010100,
20'b00010110110101100010,
20'b00010111001000110110,
20'b00010111011100010000,
20'b00010111101111110001,
20'b00011000000011011000,
20'b00011000010111000101,
20'b00011000101010111000,
20'b00011000111110110001,
20'b00011001010010110000,
20'b00011001100110110101,
20'b00011001111011000001,
20'b00011010001111010010,
20'b00011010100011101000,
20'b00011010111000000101,
20'b00011011001100100111,
20'b00011011100001010000,
20'b00011011110101111101,
20'b00011100001010110001,
20'b00011100011111101001,
20'b00011100110100101000,
20'b00011101001001101011,
20'b00011101011110110101,
20'b00011101110100000011,
20'b00011110001001010111,
20'b00011110011110110000,
20'b00011110110100001110,
20'b00011111001001110001,
20'b00011111011111011010,
20'b00011111110101000111,
20'b00100000001010111001,
20'b00100000100000110001,
20'b00100000110110101101,
20'b00100001001100101110,
20'b00100001100010110011,
20'b00100001111000111110,
20'b00100010001111001101,
20'b00100010100101100001,
20'b00100010111011111001,
20'b00100011010010010101,
20'b00100011101000110111,
20'b00100011111111011100,
20'b00100100010110000110,
20'b00100100101100110100,
20'b00100101000011100110,
20'b00100101011010011101,
20'b00100101110001011000,
20'b00100110001000010110,
20'b00100110011111011001,
20'b00100110110110011111,
20'b00100111001101101010,
20'b00100111100100111000,
20'b00100111111100001010,
20'b00101000010011100000,
20'b00101000101010111010,
20'b00101001000010010111,
20'b00101001011001110111,
20'b00101001110001011100,
20'b00101010001001000011,
20'b00101010100000101110,
20'b00101010111000011100,
20'b00101011010000001110,
20'b00101011101000000010,
20'b00101011111111111010,
20'b00101100010111110101,
20'b00101100101111110011,
20'b00101101000111110100,
20'b00101101011111111000,
20'b00101101110111111111,
20'b00101110010000001000,
20'b00101110101000010101,
20'b00101111000000100100,
20'b00101111011000110101,
20'b00101111110001001001,
20'b00110000001001100000,
20'b00110000100001111001,
20'b00110000111010010101,
20'b00110001010010110011,
20'b00110001101011010011,
20'b00110010000011110101,
20'b00110010011100011001,
20'b00110010110101000000,
20'b00110011001101101001,
20'b00110011100110010011,
20'b00110011111111000000,
20'b00110100010111101110,
20'b00110100110000011110,
20'b00110101001001010000,
20'b00110101100010000100,
20'b00110101111010111001,
20'b00110110010011110000,
20'b00110110101100101000,
20'b00110111000101100010,
20'b00110111011110011101,
20'b00110111110111011001,
20'b00111000010000010111,
20'b00111000101001010101,
20'b00111001000010010101,
20'b00111001011011010110,
20'b00111001110100011000,
20'b00111010001101011011,
20'b00111010100110011111,
20'b00111010111111100100,
20'b00111011011000101010,
20'b00111011110001110000,
20'b00111100001010110111,
20'b00111100100011111110,
20'b00111100111101000110,
20'b00111101010110001111,
20'b00111101101111011000,
20'b00111110001000100001,
20'b00111110100001101010,
20'b00111110111010110100,
20'b00111111010011111110,
20'b00111111101101001000,
20'b01000000000110010010,
20'b01000000011111011100,
20'b01000000111000100110,
20'b01000001010001110000,
20'b01000001101010111010,
20'b01000010000100000011,
20'b01000010011101001100,
20'b01000010110110010101,
20'b01000011001111011101,
20'b01000011101000100101,
20'b01000100000001101100,
20'b01000100011010110010,
20'b01000100110011111000,
20'b01000101001100111101,
20'b01000101100110000010,
20'b01000101111111000101,
20'b01000110011000001000,
20'b01000110110001001001,
20'b01000111001010001010,
20'b01000111100011001001,
20'b01000111111100000111,
20'b01001000010101000100,
20'b01001000101110000000,
20'b01001001000110111010,
20'b01001001011111110011,
20'b01001001111000101011,
20'b01001010010001100001,
20'b01001010101010010101,
20'b01001011000011001000,
20'b01001011011011111001,
20'b01001011110100101000,
20'b01001100001101010110,
20'b01001100100110000001,
20'b01001100111110101011,
20'b01001101010111010011,
20'b01001101101111111000,
20'b01001110001000011011,
20'b01001110100000111101,
20'b01001110111001011100,
20'b01001111010001111000,
20'b01001111101010010011,
20'b01010000000010101011,
20'b01010000011011000000,
20'b01010000110011010011,
20'b01010001001011100011,
20'b01010001100011110001,
20'b01010001111011111100,
20'b01010010010100000100,
20'b01010010101100001001,
20'b01010011000100001100,
20'b01010011011100001011,
20'b01010011110100001000,
20'b01010100001100000001,
20'b01010100100011110111,
20'b01010100111011101010,
20'b01010101010011011010,
20'b01010101101011000111,
20'b01010110000010110000,
20'b01010110011010010110,
20'b01010110110001111000,
20'b01010111001001010111,
20'b01010111100000110011,
20'b01010111111000001010,
20'b01011000001111011110,
20'b01011000100110101110,
20'b01011000111101111011,
20'b01011001010101000011,
20'b01011001101100001000,
20'b01011010000011001001,
20'b01011010011010000101,
20'b01011010110000111110,
20'b01011011000111110010,
20'b01011011011110100010,
20'b01011011110101001110,
20'b01011100001011110110,
20'b01011100100010011010,
20'b01011100111000111000,
20'b01011101001111010011,
20'b01011101100101101001,
20'b01011101111011111010,
20'b01011110010010000111,
20'b01011110101000001111,
20'b01011110111110010010,
20'b01011111010100010001,
20'b01011111101010001011,
20'b01011111111111111111,
20'b01100000010101101111,
20'b01100000101011011010,
20'b01100001000001000000,
20'b01100001010110100001,
20'b01100001101011111100,
20'b01100010000001010011,
20'b01100010010110100100,
20'b01100010101011110000,
20'b01100011000000110110,
20'b01100011010101110111,
20'b01100011101010110011,
20'b01100011111111101001,
20'b01100100010100011001,
20'b01100100101001000100,
20'b01100100111101101001,
20'b01100101010010001001,
20'b01100101100110100011,
20'b01100101111010110111,
20'b01100110001111000101,
20'b01100110100011001101,
20'b01100110110111001111,
20'b01100111001011001011,
20'b01100111011111000010,
20'b01100111110010110010,
20'b01101000000110011100,
20'b01101000011001111111,
20'b01101000101101011101,
20'b01101001000000110100,
20'b01101001010100000101,
20'b01101001100111001111,
20'b01101001111010010011,
20'b01101010001101010001,
20'b01101010100000001000,
20'b01101010110010111000,
20'b01101011000101100010,
20'b01101011011000000101,
20'b01101011101010100010,
20'b01101011111100111000,
20'b01101100001111000111,
20'b01101100100001001111,
20'b01101100110011010000,
20'b01101101000101001010,
20'b01101101010110111110,
20'b01101101101000101010,
20'b01101101111010001111,
20'b01101110001011101110,
20'b01101110011101000101,
20'b01101110101110010101,
20'b01101110111111011101,
20'b01101111010000011111,
20'b01101111100001011001,
20'b01101111110010001100,
20'b01110000000010110111,
20'b01110000010011011011,
20'b01110000100011110111,
20'b01110000110100001100,
20'b01110001000100011010,
20'b01110001010100100000,
20'b01110001100100011110,
20'b01110001110100010101,
20'b01110010000100000011,
20'b01110010010011101011,
20'b01110010100011001010,
20'b01110010110010100010,
20'b01110011000001110001,
20'b01110011010000111001,
20'b01110011011111111001,
20'b01110011101110110001,
20'b01110011111101100001,
20'b01110100001100001001,
20'b01110100011010101001,
20'b01110100101001000001,
20'b01110100110111010000,
20'b01110101000101011000,
20'b01110101010011010111,
20'b01110101100001001110,
20'b01110101101110111101,
20'b01110101111100100011,
20'b01110110001010000001,
20'b01110110010111010111,
20'b01110110100100100101,
20'b01110110110001101001,
20'b01110110111110100110,
20'b01110111001011011010,
20'b01110111011000000101,
20'b01110111100100101000,
20'b01110111110001000011,
20'b01110111111101010100,
20'b01111000001001011101,
20'b01111000010101011110,
20'b01111000100001010101,
20'b01111000101101000100,
20'b01111000111000101010,
20'b01111001000100001000,
20'b01111001001111011100,
20'b01111001011010101000,
20'b01111001100101101011,
20'b01111001110000100101,
20'b01111001111011010110,
20'b01111010000101111110,
20'b01111010010000011101,
20'b01111010011010110011,
20'b01111010100101000000,
20'b01111010101111000100,
20'b01111010111000111111,
20'b01111011000010110001,
20'b01111011001100011010,
20'b01111011010101111001,
20'b01111011011111010000,
20'b01111011101000011101,
20'b01111011110001100001,
20'b01111011111010011100,
20'b01111100000011001101,
20'b01111100001011110101,
20'b01111100010100010100,
20'b01111100011100101010,
20'b01111100100100110110,
20'b01111100101100111001,
20'b01111100110100110011,
20'b01111100111100100011,
20'b01111101000100001001,
20'b01111101001011100111,
20'b01111101010010111010,
20'b01111101011010000101,
20'b01111101100001000110,
20'b01111101100111111101,
20'b01111101101110101011,
20'b01111101110101001111,
20'b01111101111011101010,
20'b01111110000001111011,
20'b01111110001000000011,
20'b01111110001110000001,
20'b01111110010011110101,
20'b01111110011001100000,
20'b01111110011111000001,
20'b01111110100100011000,
20'b01111110101001100110,
20'b01111110101110101010,
20'b01111110110011100101,
20'b01111110111000010101,
20'b01111110111100111100,
20'b01111111000001011010,
20'b01111111000101101101,
20'b01111111001001110111,
20'b01111111001101110111,
20'b01111111010001101101,
20'b01111111010101011010,
20'b01111111011000111100,
20'b01111111011100010101,
20'b01111111011111100100,
20'b01111111100010101010,
20'b01111111100101100101,
20'b01111111101000010111,
20'b01111111101010111111,
20'b01111111101101011100,
20'b01111111101111110001,
20'b01111111110001111011,
20'b01111111110011111011,
20'b01111111110101110010,
20'b01111111110111011111,
20'b01111111111001000001,
20'b01111111111010011010,
20'b01111111111011101001,
20'b01111111111100101111,
20'b01111111111101101010,
20'b01111111111110011011,
20'b01111111111111000011,
20'b01111111111111100001,
20'b01111111111111110100,
20'b01111111111111111110,
20'b01111111111111111110,
20'b01111111111111110100,
20'b01111111111111100001,
20'b01111111111111000011,
20'b01111111111110011011,
20'b01111111111101101010,
20'b01111111111100101111,
20'b01111111111011101001,
20'b01111111111010011010,
20'b01111111111001000001,
20'b01111111110111011111,
20'b01111111110101110010,
20'b01111111110011111011,
20'b01111111110001111011,
20'b01111111101111110001,
20'b01111111101101011100,
20'b01111111101010111111,
20'b01111111101000010111,
20'b01111111100101100101,
20'b01111111100010101010,
20'b01111111011111100100,
20'b01111111011100010101,
20'b01111111011000111100,
20'b01111111010101011010,
20'b01111111010001101101,
20'b01111111001101110111,
20'b01111111001001110111,
20'b01111111000101101101,
20'b01111111000001011010,
20'b01111110111100111100,
20'b01111110111000010101,
20'b01111110110011100101,
20'b01111110101110101010,
20'b01111110101001100110,
20'b01111110100100011000,
20'b01111110011111000001,
20'b01111110011001100000,
20'b01111110010011110101,
20'b01111110001110000001,
20'b01111110001000000011,
20'b01111110000001111011,
20'b01111101111011101010,
20'b01111101110101001111,
20'b01111101101110101011,
20'b01111101100111111101,
20'b01111101100001000110,
20'b01111101011010000101,
20'b01111101010010111010,
20'b01111101001011100111,
20'b01111101000100001001,
20'b01111100111100100011,
20'b01111100110100110011,
20'b01111100101100111001,
20'b01111100100100110110,
20'b01111100011100101010,
20'b01111100010100010100,
20'b01111100001011110101,
20'b01111100000011001101,
20'b01111011111010011100,
20'b01111011110001100001,
20'b01111011101000011101,
20'b01111011011111010000,
20'b01111011010101111001,
20'b01111011001100011010,
20'b01111011000010110001,
20'b01111010111000111111,
20'b01111010101111000100,
20'b01111010100101000000,
20'b01111010011010110011,
20'b01111010010000011101,
20'b01111010000101111110,
20'b01111001111011010110,
20'b01111001110000100101,
20'b01111001100101101011,
20'b01111001011010101000,
20'b01111001001111011100,
20'b01111001000100001000,
20'b01111000111000101010,
20'b01111000101101000100,
20'b01111000100001010101,
20'b01111000010101011110,
20'b01111000001001011101,
20'b01110111111101010100,
20'b01110111110001000011,
20'b01110111100100101000,
20'b01110111011000000101,
20'b01110111001011011010,
20'b01110110111110100110,
20'b01110110110001101001,
20'b01110110100100100101,
20'b01110110010111010111,
20'b01110110001010000001,
20'b01110101111100100011,
20'b01110101101110111101,
20'b01110101100001001110,
20'b01110101010011010111,
20'b01110101000101011000,
20'b01110100110111010000,
20'b01110100101001000001,
20'b01110100011010101001,
20'b01110100001100001001,
20'b01110011111101100001,
20'b01110011101110110001,
20'b01110011011111111001,
20'b01110011010000111001,
20'b01110011000001110001,
20'b01110010110010100010,
20'b01110010100011001010,
20'b01110010010011101011,
20'b01110010000100000011,
20'b01110001110100010101,
20'b01110001100100011110,
20'b01110001010100100000,
20'b01110001000100011010,
20'b01110000110100001100,
20'b01110000100011110111,
20'b01110000010011011011,
20'b01110000000010110111,
20'b01101111110010001100,
20'b01101111100001011001,
20'b01101111010000011111,
20'b01101110111111011101,
20'b01101110101110010101,
20'b01101110011101000101,
20'b01101110001011101110,
20'b01101101111010001111,
20'b01101101101000101010,
20'b01101101010110111110,
20'b01101101000101001010,
20'b01101100110011010000,
20'b01101100100001001111,
20'b01101100001111000111,
20'b01101011111100111000,
20'b01101011101010100010,
20'b01101011011000000101,
20'b01101011000101100010,
20'b01101010110010111000,
20'b01101010100000001000,
20'b01101010001101010001,
20'b01101001111010010011,
20'b01101001100111001111,
20'b01101001010100000101,
20'b01101001000000110100,
20'b01101000101101011101,
20'b01101000011001111111,
20'b01101000000110011100,
20'b01100111110010110010,
20'b01100111011111000010,
20'b01100111001011001011,
20'b01100110110111001111,
20'b01100110100011001101,
20'b01100110001111000101,
20'b01100101111010110111,
20'b01100101100110100011,
20'b01100101010010001001,
20'b01100100111101101001,
20'b01100100101001000100,
20'b01100100010100011001,
20'b01100011111111101001,
20'b01100011101010110011,
20'b01100011010101110111,
20'b01100011000000110110,
20'b01100010101011110000,
20'b01100010010110100100,
20'b01100010000001010011,
20'b01100001101011111100,
20'b01100001010110100001,
20'b01100001000001000000,
20'b01100000101011011010,
20'b01100000010101101111,
20'b01100000000000000000,
20'b01011111101010001011,
20'b01011111010100010001,
20'b01011110111110010010,
20'b01011110101000001111,
20'b01011110010010000111,
20'b01011101111011111010,
20'b01011101100101101001,
20'b01011101001111010011,
20'b01011100111000111000,
20'b01011100100010011010,
20'b01011100001011110110,
20'b01011011110101001110,
20'b01011011011110100010,
20'b01011011000111110010,
20'b01011010110000111110,
20'b01011010011010000101,
20'b01011010000011001001,
20'b01011001101100001000,
20'b01011001010101000011,
20'b01011000111101111011,
20'b01011000100110101110,
20'b01011000001111011110,
20'b01010111111000001010,
20'b01010111100000110011,
20'b01010111001001010111,
20'b01010110110001111000,
20'b01010110011010010110,
20'b01010110000010110000,
20'b01010101101011000111,
20'b01010101010011011010,
20'b01010100111011101010,
20'b01010100100011110111,
20'b01010100001100000001,
20'b01010011110100001000,
20'b01010011011100001011,
20'b01010011000100001100,
20'b01010010101100001001,
20'b01010010010100000100,
20'b01010001111011111100,
20'b01010001100011110001,
20'b01010001001011100011,
20'b01010000110011010011,
20'b01010000011011000000,
20'b01010000000010101011,
20'b01001111101010010011,
20'b01001111010001111000,
20'b01001110111001011100,
20'b01001110100000111101,
20'b01001110001000011011,
20'b01001101101111111000,
20'b01001101010111010011,
20'b01001100111110101011,
20'b01001100100110000001,
20'b01001100001101010110,
20'b01001011110100101000,
20'b01001011011011111001,
20'b01001011000011001000,
20'b01001010101010010101,
20'b01001010010001100001,
20'b01001001111000101011,
20'b01001001011111110011,
20'b01001001000110111010,
20'b01001000101110000000,
20'b01001000010101000100,
20'b01000111111100000111,
20'b01000111100011001001,
20'b01000111001010001010,
20'b01000110110001001001,
20'b01000110011000001000,
20'b01000101111111000101,
20'b01000101100110000010,
20'b01000101001100111101,
20'b01000100110011111000,
20'b01000100011010110010,
20'b01000100000001101100,
20'b01000011101000100101,
20'b01000011001111011101,
20'b01000010110110010101,
20'b01000010011101001100,
20'b01000010000100000011,
20'b01000001101010111010,
20'b01000001010001110000,
20'b01000000111000100110,
20'b01000000011111011100,
20'b01000000000110010010,
20'b00111111101101001000,
20'b00111111010011111110,
20'b00111110111010110100,
20'b00111110100001101010,
20'b00111110001000100001,
20'b00111101101111011000,
20'b00111101010110001111,
20'b00111100111101000110,
20'b00111100100011111110,
20'b00111100001010110111,
20'b00111011110001110000,
20'b00111011011000101010,
20'b00111010111111100100,
20'b00111010100110011111,
20'b00111010001101011011,
20'b00111001110100011000,
20'b00111001011011010110,
20'b00111001000010010101,
20'b00111000101001010101,
20'b00111000010000010111,
20'b00110111110111011001,
20'b00110111011110011101,
20'b00110111000101100010,
20'b00110110101100101000,
20'b00110110010011110000,
20'b00110101111010111001,
20'b00110101100010000100,
20'b00110101001001010000,
20'b00110100110000011110,
20'b00110100010111101110,
20'b00110011111111000000,
20'b00110011100110010011,
20'b00110011001101101001,
20'b00110010110101000000,
20'b00110010011100011001,
20'b00110010000011110101,
20'b00110001101011010011,
20'b00110001010010110011,
20'b00110000111010010101,
20'b00110000100001111001,
20'b00110000001001100000,
20'b00101111110001001001,
20'b00101111011000110101,
20'b00101111000000100100,
20'b00101110101000010101,
20'b00101110010000001000,
20'b00101101110111111111,
20'b00101101011111111000,
20'b00101101000111110100,
20'b00101100101111110011,
20'b00101100010111110101,
20'b00101011111111111010,
20'b00101011101000000010,
20'b00101011010000001110,
20'b00101010111000011100,
20'b00101010100000101110,
20'b00101010001001000011,
20'b00101001110001011100,
20'b00101001011001110111,
20'b00101001000010010111,
20'b00101000101010111010,
20'b00101000010011100000,
20'b00100111111100001010,
20'b00100111100100111000,
20'b00100111001101101010,
20'b00100110110110011111,
20'b00100110011111011001,
20'b00100110001000010110,
20'b00100101110001011000,
20'b00100101011010011101,
20'b00100101000011100110,
20'b00100100101100110100,
20'b00100100010110000110,
20'b00100011111111011100,
20'b00100011101000110111,
20'b00100011010010010101,
20'b00100010111011111001,
20'b00100010100101100001,
20'b00100010001111001101,
20'b00100001111000111110,
20'b00100001100010110011,
20'b00100001001100101110,
20'b00100000110110101101,
20'b00100000100000110001,
20'b00100000001010111001,
20'b00011111110101000111,
20'b00011111011111011010,
20'b00011111001001110001,
20'b00011110110100001110,
20'b00011110011110110000,
20'b00011110001001010111,
20'b00011101110100000011,
20'b00011101011110110101,
20'b00011101001001101011,
20'b00011100110100101000,
20'b00011100011111101001,
20'b00011100001010110001,
20'b00011011110101111101,
20'b00011011100001010000,
20'b00011011001100100111,
20'b00011010111000000101,
20'b00011010100011101000,
20'b00011010001111010010,
20'b00011001111011000001,
20'b00011001100110110101,
20'b00011001010010110000,
20'b00011000111110110001,
20'b00011000101010111000,
20'b00011000010111000101,
20'b00011000000011011000,
20'b00010111101111110001,
20'b00010111011100010000,
20'b00010111001000110110,
20'b00010110110101100010,
20'b00010110100010010100,
20'b00010110001111001101,
20'b00010101111100001100,
20'b00010101101001010010,
20'b00010101010110011110,
20'b00010101000011110001,
20'b00010100110001001010,
20'b00010100011110101010,
20'b00010100001100010001,
20'b00010011111001111111,
20'b00010011100111110011,
20'b00010011010101101111,
20'b00010011000011110001,
20'b00010010110001111010,
20'b00010010100000001010,
20'b00010010001110100001,
20'b00010001111101000000,
20'b00010001101011100101,
20'b00010001011010010001,
20'b00010001001001000101,
20'b00010000111000000000,
20'b00010000100111000010,
20'b00010000010110001100,
20'b00010000000101011101,
20'b00001111110100110101,
20'b00001111100100010101,
20'b00001111010011111100,
20'b00001111000011101011,
20'b00001110110011100001,
20'b00001110100011011111,
20'b00001110010011100101,
20'b00001110000011110010,
20'b00001101110100000111,
20'b00001101100100100100,
20'b00001101010101001000,
20'b00001101000101110101,
20'b00001100110110101001,
20'b00001100100111100101,
20'b00001100011000101001,
20'b00001100001001110101,
20'b00001011111011001001,
20'b00001011101100100101,
20'b00001011011110001001,
20'b00001011001111110110,
20'b00001011000001101010,
20'b00001010110011100111,
20'b00001010100101101011,
20'b00001010010111111001,
20'b00001010001010001110,
20'b00001001111100101100,
20'b00001001101111010010,
20'b00001001100010000000,
20'b00001001010100110111,
20'b00001001000111110110,
20'b00001000111010111110,
20'b00001000101110001110,
20'b00001000100001100111,
20'b00001000010101001001,
20'b00001000001000110011,
20'b00000111111100100101,
20'b00000111110000100000,
20'b00000111100100100100,
20'b00000111011000110001,
20'b00000111001101000111,
20'b00000111000001100101,
20'b00000110110110001100,
20'b00000110101010111100,
20'b00000110011111110100,
20'b00000110010100110110,
20'b00000110001010000001,
20'b00000101111111010100,
20'b00000101110100110000,
20'b00000101101010010110,
20'b00000101100000000100,
20'b00000101010101111100,
20'b00000101001011111100,
20'b00000101000010000110,
20'b00000100111000011001,
20'b00000100101110110100,
20'b00000100100101011001,
20'b00000100011100001000,
20'b00000100010010111111,
20'b00000100001010000000,
20'b00000100000001001001,
20'b00000011111000011101,
20'b00000011101111111001,
20'b00000011100111011111,
20'b00000011011111001110,
20'b00000011010111000110,
20'b00000011001111001000,
20'b00000011000111010011,
20'b00000010111111101000,
20'b00000010111000000110,
20'b00000010110000101101,
20'b00000010101001011110,
20'b00000010100010011001,
20'b00000010011011011100,
20'b00000010010100101010,
20'b00000010001110000001,
20'b00000010000111100001,
20'b00000010000001001011,
20'b00000001111010111111,
20'b00000001110100111100,
20'b00000001101111000011,
20'b00000001101001010011,
20'b00000001100011101101,
20'b00000001011110010001,
20'b00000001011000111111,
20'b00000001010011110110,
20'b00000001001110110110,
20'b00000001001010000001,
20'b00000001000101010101,
20'b00000001000000110011,
20'b00000000111100011010,
20'b00000000111000001100,
20'b00000000110100000111,
20'b00000000110000001100,
20'b00000000101100011010,
20'b00000000101000110011,
20'b00000000100101010101,
20'b00000000100010000001,
20'b00000000011110110111,
20'b00000000011011110110,
20'b00000000011001000000,
20'b00000000010110010011,
20'b00000000010011110000,
20'b00000000010001010111,
20'b00000000001111001000,
20'b00000000001101000011,
20'b00000000001011000111,
20'b00000000001001010110,
20'b00000000000111101110,
20'b00000000000110010000,
20'b00000000000100111100,
20'b00000000000011110010,
20'b00000000000010110001,
20'b00000000000001111011,
20'b00000000000001001111,
20'b00000000000000101100,
20'b00000000000000010011,
20'b00000000000000000100,
20'b00000000000000000000
};

`endif