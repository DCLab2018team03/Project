`ifndef _ACAPPELLA_DEFINE_VH_
`define _ACAPPELLA_DEFINE_VH_

// TODO
// Divide the SDRAM into reasonable chunks