`ifndef _ACAPPELLA_DEFINE_SV_
`define _ACAPPELLA_DEFINE_SV_

// TODO
// Divide the SDRAM into reasonable chunks

paramater WindowSize = 512; // window size for time-stretching and pitch-shifting
