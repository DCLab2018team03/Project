`ifndef _PITCH_DEFINE_SV_
`define _PITCH_DEFINE_SV_
// window size for time-stretching and pitch-shifting, if you change the window size,
// remember to modify the hanning coefficients below
parameter WindowSize = 512; 

// hanning window parameter 0~512
// format: unsigned, the first bit is preserverd (in case they are used to be signed),
//         the remaining represents the floating point of the coefficients
//         (no precise 1 occurs, so it's OK not to store the int part)
parameter [15:0] HANN_C000 = 16'b0000000000000000;
parameter [15:0] HANN_C001 = 16'b0000000000000001;
parameter [15:0] HANN_C002 = 16'b0000000000000100;
parameter [15:0] HANN_C003 = 16'b0000000000001011;
parameter [15:0] HANN_C004 = 16'b0000000000010011;
parameter [15:0] HANN_C005 = 16'b0000000000011110;
parameter [15:0] HANN_C006 = 16'b0000000000101100;
parameter [15:0] HANN_C007 = 16'b0000000000111100;
parameter [15:0] HANN_C008 = 16'b0000000001001111;
parameter [15:0] HANN_C009 = 16'b0000000001100100;
parameter [15:0] HANN_C010 = 16'b0000000001111011;
parameter [15:0] HANN_C011 = 16'b0000000010010101;
parameter [15:0] HANN_C012 = 16'b0000000010110010;
parameter [15:0] HANN_C013 = 16'b0000000011010000;
parameter [15:0] HANN_C014 = 16'b0000000011110010;
parameter [15:0] HANN_C015 = 16'b0000000100010101;
parameter [15:0] HANN_C016 = 16'b0000000100111100;
parameter [15:0] HANN_C017 = 16'b0000000101100100;
parameter [15:0] HANN_C018 = 16'b0000000110001111;
parameter [15:0] HANN_C019 = 16'b0000000110111101;
parameter [15:0] HANN_C020 = 16'b0000000111101100;
parameter [15:0] HANN_C021 = 16'b0000001000011111;
parameter [15:0] HANN_C022 = 16'b0000001001010011;
parameter [15:0] HANN_C023 = 16'b0000001010001010;
parameter [15:0] HANN_C024 = 16'b0000001011000100;
parameter [15:0] HANN_C025 = 16'b0000001100000000;
parameter [15:0] HANN_C026 = 16'b0000001100111110;
parameter [15:0] HANN_C027 = 16'b0000001101111110;
parameter [15:0] HANN_C028 = 16'b0000001111000001;
parameter [15:0] HANN_C029 = 16'b0000010000000110;
parameter [15:0] HANN_C030 = 16'b0000010001001110;
parameter [15:0] HANN_C031 = 16'b0000010010010111;
parameter [15:0] HANN_C032 = 16'b0000010011100011;
parameter [15:0] HANN_C033 = 16'b0000010100110010;
parameter [15:0] HANN_C034 = 16'b0000010110000011;
parameter [15:0] HANN_C035 = 16'b0000010111010101;
parameter [15:0] HANN_C036 = 16'b0000011000101011;
parameter [15:0] HANN_C037 = 16'b0000011010000010;
parameter [15:0] HANN_C038 = 16'b0000011011011100;
parameter [15:0] HANN_C039 = 16'b0000011100110111;
parameter [15:0] HANN_C040 = 16'b0000011110010110;
parameter [15:0] HANN_C041 = 16'b0000011111110110;
parameter [15:0] HANN_C042 = 16'b0000100001011000;
parameter [15:0] HANN_C043 = 16'b0000100010111101;
parameter [15:0] HANN_C044 = 16'b0000100100100011;
parameter [15:0] HANN_C045 = 16'b0000100110001100;
parameter [15:0] HANN_C046 = 16'b0000100111110111;
parameter [15:0] HANN_C047 = 16'b0000101001100100;
parameter [15:0] HANN_C048 = 16'b0000101011010011;
parameter [15:0] HANN_C049 = 16'b0000101101000100;
parameter [15:0] HANN_C050 = 16'b0000101110111000;
parameter [15:0] HANN_C051 = 16'b0000110000101101;
parameter [15:0] HANN_C052 = 16'b0000110010100100;
parameter [15:0] HANN_C053 = 16'b0000110100011101;
parameter [15:0] HANN_C054 = 16'b0000110110011000;
parameter [15:0] HANN_C055 = 16'b0000111000010101;
parameter [15:0] HANN_C056 = 16'b0000111010010100;
parameter [15:0] HANN_C057 = 16'b0000111100010101;
parameter [15:0] HANN_C058 = 16'b0000111110011000;
parameter [15:0] HANN_C059 = 16'b0001000000011101;
parameter [15:0] HANN_C060 = 16'b0001000010100100;
parameter [15:0] HANN_C061 = 16'b0001000100101100;
parameter [15:0] HANN_C062 = 16'b0001000110110110;
parameter [15:0] HANN_C063 = 16'b0001001001000010;
parameter [15:0] HANN_C064 = 16'b0001001011010000;
parameter [15:0] HANN_C065 = 16'b0001001101100000;
parameter [15:0] HANN_C066 = 16'b0001001111110001;
parameter [15:0] HANN_C067 = 16'b0001010010000100;
parameter [15:0] HANN_C068 = 16'b0001010100011001;
parameter [15:0] HANN_C069 = 16'b0001010110101111;
parameter [15:0] HANN_C070 = 16'b0001011001000111;
parameter [15:0] HANN_C071 = 16'b0001011011100000;
parameter [15:0] HANN_C072 = 16'b0001011101111100;
parameter [15:0] HANN_C073 = 16'b0001100000011000;
parameter [15:0] HANN_C074 = 16'b0001100010110111;
parameter [15:0] HANN_C075 = 16'b0001100101010110;
parameter [15:0] HANN_C076 = 16'b0001100111111000;
parameter [15:0] HANN_C077 = 16'b0001101010011010;
parameter [15:0] HANN_C078 = 16'b0001101100111111;
parameter [15:0] HANN_C079 = 16'b0001101111100100;
parameter [15:0] HANN_C080 = 16'b0001110010001011;
parameter [15:0] HANN_C081 = 16'b0001110100110100;
parameter [15:0] HANN_C082 = 16'b0001110111011101;
parameter [15:0] HANN_C083 = 16'b0001111010001000;
parameter [15:0] HANN_C084 = 16'b0001111100110101;
parameter [15:0] HANN_C085 = 16'b0001111111100010;
parameter [15:0] HANN_C086 = 16'b0010000010010001;
parameter [15:0] HANN_C087 = 16'b0010000101000001;
parameter [15:0] HANN_C088 = 16'b0010000111110011;
parameter [15:0] HANN_C089 = 16'b0010001010100101;
parameter [15:0] HANN_C090 = 16'b0010001101011001;
parameter [15:0] HANN_C091 = 16'b0010010000001101;
parameter [15:0] HANN_C092 = 16'b0010010011000011;
parameter [15:0] HANN_C093 = 16'b0010010101111010;
parameter [15:0] HANN_C094 = 16'b0010011000110010;
parameter [15:0] HANN_C095 = 16'b0010011011101011;
parameter [15:0] HANN_C096 = 16'b0010011110100101;
parameter [15:0] HANN_C097 = 16'b0010100001011111;
parameter [15:0] HANN_C098 = 16'b0010100100011011;
parameter [15:0] HANN_C099 = 16'b0010100111011000;
parameter [15:0] HANN_C100 = 16'b0010101010010101;
parameter [15:0] HANN_C101 = 16'b0010101101010011;
parameter [15:0] HANN_C102 = 16'b0010110000010010;
parameter [15:0] HANN_C103 = 16'b0010110011010010;
parameter [15:0] HANN_C104 = 16'b0010110110010011;
parameter [15:0] HANN_C105 = 16'b0010111001010100;
parameter [15:0] HANN_C106 = 16'b0010111100010110;
parameter [15:0] HANN_C107 = 16'b0010111111011001;
parameter [15:0] HANN_C108 = 16'b0011000010011100;
parameter [15:0] HANN_C109 = 16'b0011000101100000;
parameter [15:0] HANN_C110 = 16'b0011001000100100;
parameter [15:0] HANN_C111 = 16'b0011001011101001;
parameter [15:0] HANN_C112 = 16'b0011001110101110;
parameter [15:0] HANN_C113 = 16'b0011010001110100;
parameter [15:0] HANN_C114 = 16'b0011010100111011;
parameter [15:0] HANN_C115 = 16'b0011011000000001;
parameter [15:0] HANN_C116 = 16'b0011011011001001;
parameter [15:0] HANN_C117 = 16'b0011011110010000;
parameter [15:0] HANN_C118 = 16'b0011100001011000;
parameter [15:0] HANN_C119 = 16'b0011100100100000;
parameter [15:0] HANN_C120 = 16'b0011100111101001;
parameter [15:0] HANN_C121 = 16'b0011101010110001;
parameter [15:0] HANN_C122 = 16'b0011101101111010;
parameter [15:0] HANN_C123 = 16'b0011110001000011;
parameter [15:0] HANN_C124 = 16'b0011110100001100;
parameter [15:0] HANN_C125 = 16'b0011110111010110;
parameter [15:0] HANN_C126 = 16'b0011111010011111;
parameter [15:0] HANN_C127 = 16'b0011111101101000;
parameter [15:0] HANN_C128 = 16'b0100000000110010;
parameter [15:0] HANN_C129 = 16'b0100000011111011;
parameter [15:0] HANN_C130 = 16'b0100000111000101;
parameter [15:0] HANN_C131 = 16'b0100001010001110;
parameter [15:0] HANN_C132 = 16'b0100001101010111;
parameter [15:0] HANN_C133 = 16'b0100010000100000;
parameter [15:0] HANN_C134 = 16'b0100010011101001;
parameter [15:0] HANN_C135 = 16'b0100010110110010;
parameter [15:0] HANN_C136 = 16'b0100011001111011;
parameter [15:0] HANN_C137 = 16'b0100011101000011;
parameter [15:0] HANN_C138 = 16'b0100100000001011;
parameter [15:0] HANN_C139 = 16'b0100100011010011;
parameter [15:0] HANN_C140 = 16'b0100100110011010;
parameter [15:0] HANN_C141 = 16'b0100101001100001;
parameter [15:0] HANN_C142 = 16'b0100101100101000;
parameter [15:0] HANN_C143 = 16'b0100101111101110;
parameter [15:0] HANN_C144 = 16'b0100110010110011;
parameter [15:0] HANN_C145 = 16'b0100110101111001;
parameter [15:0] HANN_C146 = 16'b0100111000111101;
parameter [15:0] HANN_C147 = 16'b0100111100000001;
parameter [15:0] HANN_C148 = 16'b0100111111000101;
parameter [15:0] HANN_C149 = 16'b0101000010001000;
parameter [15:0] HANN_C150 = 16'b0101000101001010;
parameter [15:0] HANN_C151 = 16'b0101001000001100;
parameter [15:0] HANN_C152 = 16'b0101001011001101;
parameter [15:0] HANN_C153 = 16'b0101001110001101;
parameter [15:0] HANN_C154 = 16'b0101010001001100;
parameter [15:0] HANN_C155 = 16'b0101010100001011;
parameter [15:0] HANN_C156 = 16'b0101010111001001;
parameter [15:0] HANN_C157 = 16'b0101011010000110;
parameter [15:0] HANN_C158 = 16'b0101011101000010;
parameter [15:0] HANN_C159 = 16'b0101011111111101;
parameter [15:0] HANN_C160 = 16'b0101100010111000;
parameter [15:0] HANN_C161 = 16'b0101100101110001;
parameter [15:0] HANN_C162 = 16'b0101101000101001;
parameter [15:0] HANN_C163 = 16'b0101101011100001;
parameter [15:0] HANN_C164 = 16'b0101101110010111;
parameter [15:0] HANN_C165 = 16'b0101110001001100;
parameter [15:0] HANN_C166 = 16'b0101110100000000;
parameter [15:0] HANN_C167 = 16'b0101110110110011;
parameter [15:0] HANN_C168 = 16'b0101111001100101;
parameter [15:0] HANN_C169 = 16'b0101111100010110;
parameter [15:0] HANN_C170 = 16'b0101111111000101;
parameter [15:0] HANN_C171 = 16'b0110000001110100;
parameter [15:0] HANN_C172 = 16'b0110000100100001;
parameter [15:0] HANN_C173 = 16'b0110000111001100;
parameter [15:0] HANN_C174 = 16'b0110001001110111;
parameter [15:0] HANN_C175 = 16'b0110001100100000;
parameter [15:0] HANN_C176 = 16'b0110001111000111;
parameter [15:0] HANN_C177 = 16'b0110010001101110;
parameter [15:0] HANN_C178 = 16'b0110010100010011;
parameter [15:0] HANN_C179 = 16'b0110010110110110;
parameter [15:0] HANN_C180 = 16'b0110011001011000;
parameter [15:0] HANN_C181 = 16'b0110011011111001;
parameter [15:0] HANN_C182 = 16'b0110011110011000;
parameter [15:0] HANN_C183 = 16'b0110100000110101;
parameter [15:0] HANN_C184 = 16'b0110100011010001;
parameter [15:0] HANN_C185 = 16'b0110100101101100;
parameter [15:0] HANN_C186 = 16'b0110101000000100;
parameter [15:0] HANN_C187 = 16'b0110101010011100;
parameter [15:0] HANN_C188 = 16'b0110101100110001;
parameter [15:0] HANN_C189 = 16'b0110101111000101;
parameter [15:0] HANN_C190 = 16'b0110110001010111;
parameter [15:0] HANN_C191 = 16'b0110110011100111;
parameter [15:0] HANN_C192 = 16'b0110110101110110;
parameter [15:0] HANN_C193 = 16'b0110111000000011;
parameter [15:0] HANN_C194 = 16'b0110111010001110;
parameter [15:0] HANN_C195 = 16'b0110111100010111;
parameter [15:0] HANN_C196 = 16'b0110111110011111;
parameter [15:0] HANN_C197 = 16'b0111000000100101;
parameter [15:0] HANN_C198 = 16'b0111000010101000;
parameter [15:0] HANN_C199 = 16'b0111000100101010;
parameter [15:0] HANN_C200 = 16'b0111000110101010;
parameter [15:0] HANN_C201 = 16'b0111001000101000;
parameter [15:0] HANN_C202 = 16'b0111001010100101;
parameter [15:0] HANN_C203 = 16'b0111001100011111;
parameter [15:0] HANN_C204 = 16'b0111001110010111;
parameter [15:0] HANN_C205 = 16'b0111010000001101;
parameter [15:0] HANN_C206 = 16'b0111010010000001;
parameter [15:0] HANN_C207 = 16'b0111010011110011;
parameter [15:0] HANN_C208 = 16'b0111010101100100;
parameter [15:0] HANN_C209 = 16'b0111010111010010;
parameter [15:0] HANN_C210 = 16'b0111011000111110;
parameter [15:0] HANN_C211 = 16'b0111011010100111;
parameter [15:0] HANN_C212 = 16'b0111011100001111;
parameter [15:0] HANN_C213 = 16'b0111011101110101;
parameter [15:0] HANN_C214 = 16'b0111011111011000;
parameter [15:0] HANN_C215 = 16'b0111100000111010;
parameter [15:0] HANN_C216 = 16'b0111100010011001;
parameter [15:0] HANN_C217 = 16'b0111100011110110;
parameter [15:0] HANN_C218 = 16'b0111100101010000;
parameter [15:0] HANN_C219 = 16'b0111100110101001;
parameter [15:0] HANN_C220 = 16'b0111100111111111;
parameter [15:0] HANN_C221 = 16'b0111101001010011;
parameter [15:0] HANN_C222 = 16'b0111101010100101;
parameter [15:0] HANN_C223 = 16'b0111101011110101;
parameter [15:0] HANN_C224 = 16'b0111101101000010;
parameter [15:0] HANN_C225 = 16'b0111101110001101;
parameter [15:0] HANN_C226 = 16'b0111101111010101;
parameter [15:0] HANN_C227 = 16'b0111110000011100;
parameter [15:0] HANN_C228 = 16'b0111110001100000;
parameter [15:0] HANN_C229 = 16'b0111110010100001;
parameter [15:0] HANN_C230 = 16'b0111110011100001;
parameter [15:0] HANN_C231 = 16'b0111110100011110;
parameter [15:0] HANN_C232 = 16'b0111110101011000;
parameter [15:0] HANN_C233 = 16'b0111110110010000;
parameter [15:0] HANN_C234 = 16'b0111110111000110;
parameter [15:0] HANN_C235 = 16'b0111110111111010;
parameter [15:0] HANN_C236 = 16'b0111111000101011;
parameter [15:0] HANN_C237 = 16'b0111111001011001;
parameter [15:0] HANN_C238 = 16'b0111111010000110;
parameter [15:0] HANN_C239 = 16'b0111111010101111;
parameter [15:0] HANN_C240 = 16'b0111111011010111;
parameter [15:0] HANN_C241 = 16'b0111111011111100;
parameter [15:0] HANN_C242 = 16'b0111111100011110;
parameter [15:0] HANN_C243 = 16'b0111111100111110;
parameter [15:0] HANN_C244 = 16'b0111111101011100;
parameter [15:0] HANN_C245 = 16'b0111111101110111;
parameter [15:0] HANN_C246 = 16'b0111111110010000;
parameter [15:0] HANN_C247 = 16'b0111111110100110;
parameter [15:0] HANN_C248 = 16'b0111111110111010;
parameter [15:0] HANN_C249 = 16'b0111111111001011;
parameter [15:0] HANN_C250 = 16'b0111111111011010;
parameter [15:0] HANN_C251 = 16'b0111111111100110;
parameter [15:0] HANN_C252 = 16'b0111111111110000;
parameter [15:0] HANN_C253 = 16'b0111111111111000;
parameter [15:0] HANN_C254 = 16'b0111111111111101;
parameter [15:0] HANN_C255 = 16'b0111111111111111;
// -------------------------------------------------- symmetric from here
parameter [15:0] HANN_C256 = 16'b0111111111111111;
parameter [15:0] HANN_C257 = 16'b0111111111111101;
parameter [15:0] HANN_C258 = 16'b0111111111111000;
parameter [15:0] HANN_C259 = 16'b0111111111110000;
parameter [15:0] HANN_C260 = 16'b0111111111100110;
parameter [15:0] HANN_C261 = 16'b0111111111011010;
parameter [15:0] HANN_C262 = 16'b0111111111001011;
parameter [15:0] HANN_C263 = 16'b0111111110111010;
parameter [15:0] HANN_C264 = 16'b0111111110100110;
parameter [15:0] HANN_C265 = 16'b0111111110010000;
parameter [15:0] HANN_C266 = 16'b0111111101110111;
parameter [15:0] HANN_C267 = 16'b0111111101011100;
parameter [15:0] HANN_C268 = 16'b0111111100111110;
parameter [15:0] HANN_C269 = 16'b0111111100011110;
parameter [15:0] HANN_C270 = 16'b0111111011111100;
parameter [15:0] HANN_C271 = 16'b0111111011010111;
parameter [15:0] HANN_C272 = 16'b0111111010101111;
parameter [15:0] HANN_C273 = 16'b0111111010000110;
parameter [15:0] HANN_C274 = 16'b0111111001011001;
parameter [15:0] HANN_C275 = 16'b0111111000101011;
parameter [15:0] HANN_C276 = 16'b0111110111111010;
parameter [15:0] HANN_C277 = 16'b0111110111000110;
parameter [15:0] HANN_C278 = 16'b0111110110010000;
parameter [15:0] HANN_C279 = 16'b0111110101011000;
parameter [15:0] HANN_C280 = 16'b0111110100011110;
parameter [15:0] HANN_C281 = 16'b0111110011100001;
parameter [15:0] HANN_C282 = 16'b0111110010100001;
parameter [15:0] HANN_C283 = 16'b0111110001100000;
parameter [15:0] HANN_C284 = 16'b0111110000011100;
parameter [15:0] HANN_C285 = 16'b0111101111010101;
parameter [15:0] HANN_C286 = 16'b0111101110001101;
parameter [15:0] HANN_C287 = 16'b0111101101000010;
parameter [15:0] HANN_C288 = 16'b0111101011110101;
parameter [15:0] HANN_C289 = 16'b0111101010100101;
parameter [15:0] HANN_C290 = 16'b0111101001010011;
parameter [15:0] HANN_C291 = 16'b0111100111111111;
parameter [15:0] HANN_C292 = 16'b0111100110101001;
parameter [15:0] HANN_C293 = 16'b0111100101010000;
parameter [15:0] HANN_C294 = 16'b0111100011110110;
parameter [15:0] HANN_C295 = 16'b0111100010011001;
parameter [15:0] HANN_C296 = 16'b0111100000111010;
parameter [15:0] HANN_C297 = 16'b0111011111011000;
parameter [15:0] HANN_C298 = 16'b0111011101110101;
parameter [15:0] HANN_C299 = 16'b0111011100001111;
parameter [15:0] HANN_C300 = 16'b0111011010100111;
parameter [15:0] HANN_C301 = 16'b0111011000111110;
parameter [15:0] HANN_C302 = 16'b0111010111010010;
parameter [15:0] HANN_C303 = 16'b0111010101100100;
parameter [15:0] HANN_C304 = 16'b0111010011110011;
parameter [15:0] HANN_C305 = 16'b0111010010000001;
parameter [15:0] HANN_C306 = 16'b0111010000001101;
parameter [15:0] HANN_C307 = 16'b0111001110010111;
parameter [15:0] HANN_C308 = 16'b0111001100011111;
parameter [15:0] HANN_C309 = 16'b0111001010100101;
parameter [15:0] HANN_C310 = 16'b0111001000101000;
parameter [15:0] HANN_C311 = 16'b0111000110101010;
parameter [15:0] HANN_C312 = 16'b0111000100101010;
parameter [15:0] HANN_C313 = 16'b0111000010101000;
parameter [15:0] HANN_C314 = 16'b0111000000100101;
parameter [15:0] HANN_C315 = 16'b0110111110011111;
parameter [15:0] HANN_C316 = 16'b0110111100010111;
parameter [15:0] HANN_C317 = 16'b0110111010001110;
parameter [15:0] HANN_C318 = 16'b0110111000000011;
parameter [15:0] HANN_C319 = 16'b0110110101110110;
parameter [15:0] HANN_C320 = 16'b0110110011100111;
parameter [15:0] HANN_C321 = 16'b0110110001010111;
parameter [15:0] HANN_C322 = 16'b0110101111000101;
parameter [15:0] HANN_C323 = 16'b0110101100110001;
parameter [15:0] HANN_C324 = 16'b0110101010011100;
parameter [15:0] HANN_C325 = 16'b0110101000000100;
parameter [15:0] HANN_C326 = 16'b0110100101101100;
parameter [15:0] HANN_C327 = 16'b0110100011010001;
parameter [15:0] HANN_C328 = 16'b0110100000110101;
parameter [15:0] HANN_C329 = 16'b0110011110011000;
parameter [15:0] HANN_C330 = 16'b0110011011111001;
parameter [15:0] HANN_C331 = 16'b0110011001011000;
parameter [15:0] HANN_C332 = 16'b0110010110110110;
parameter [15:0] HANN_C333 = 16'b0110010100010011;
parameter [15:0] HANN_C334 = 16'b0110010001101110;
parameter [15:0] HANN_C335 = 16'b0110001111000111;
parameter [15:0] HANN_C336 = 16'b0110001100100000;
parameter [15:0] HANN_C337 = 16'b0110001001110111;
parameter [15:0] HANN_C338 = 16'b0110000111001100;
parameter [15:0] HANN_C339 = 16'b0110000100100001;
parameter [15:0] HANN_C340 = 16'b0110000001110100;
parameter [15:0] HANN_C341 = 16'b0101111111000101;
parameter [15:0] HANN_C342 = 16'b0101111100010110;
parameter [15:0] HANN_C343 = 16'b0101111001100101;
parameter [15:0] HANN_C344 = 16'b0101110110110011;
parameter [15:0] HANN_C345 = 16'b0101110100000000;
parameter [15:0] HANN_C346 = 16'b0101110001001100;
parameter [15:0] HANN_C347 = 16'b0101101110010111;
parameter [15:0] HANN_C348 = 16'b0101101011100001;
parameter [15:0] HANN_C349 = 16'b0101101000101001;
parameter [15:0] HANN_C350 = 16'b0101100101110001;
parameter [15:0] HANN_C351 = 16'b0101100010111000;
parameter [15:0] HANN_C352 = 16'b0101011111111101;
parameter [15:0] HANN_C353 = 16'b0101011101000010;
parameter [15:0] HANN_C354 = 16'b0101011010000110;
parameter [15:0] HANN_C355 = 16'b0101010111001001;
parameter [15:0] HANN_C356 = 16'b0101010100001011;
parameter [15:0] HANN_C357 = 16'b0101010001001100;
parameter [15:0] HANN_C358 = 16'b0101001110001101;
parameter [15:0] HANN_C359 = 16'b0101001011001101;
parameter [15:0] HANN_C360 = 16'b0101001000001100;
parameter [15:0] HANN_C361 = 16'b0101000101001010;
parameter [15:0] HANN_C362 = 16'b0101000010001000;
parameter [15:0] HANN_C363 = 16'b0100111111000101;
parameter [15:0] HANN_C364 = 16'b0100111100000001;
parameter [15:0] HANN_C365 = 16'b0100111000111101;
parameter [15:0] HANN_C366 = 16'b0100110101111001;
parameter [15:0] HANN_C367 = 16'b0100110010110011;
parameter [15:0] HANN_C368 = 16'b0100101111101110;
parameter [15:0] HANN_C369 = 16'b0100101100101000;
parameter [15:0] HANN_C370 = 16'b0100101001100001;
parameter [15:0] HANN_C371 = 16'b0100100110011010;
parameter [15:0] HANN_C372 = 16'b0100100011010011;
parameter [15:0] HANN_C373 = 16'b0100100000001011;
parameter [15:0] HANN_C374 = 16'b0100011101000011;
parameter [15:0] HANN_C375 = 16'b0100011001111011;
parameter [15:0] HANN_C376 = 16'b0100010110110010;
parameter [15:0] HANN_C377 = 16'b0100010011101001;
parameter [15:0] HANN_C378 = 16'b0100010000100000;
parameter [15:0] HANN_C379 = 16'b0100001101010111;
parameter [15:0] HANN_C380 = 16'b0100001010001110;
parameter [15:0] HANN_C381 = 16'b0100000111000101;
parameter [15:0] HANN_C382 = 16'b0100000011111011;
parameter [15:0] HANN_C383 = 16'b0100000000110010;
parameter [15:0] HANN_C384 = 16'b0011111101101000;
parameter [15:0] HANN_C385 = 16'b0011111010011111;
parameter [15:0] HANN_C386 = 16'b0011110111010110;
parameter [15:0] HANN_C387 = 16'b0011110100001100;
parameter [15:0] HANN_C388 = 16'b0011110001000011;
parameter [15:0] HANN_C389 = 16'b0011101101111010;
parameter [15:0] HANN_C390 = 16'b0011101010110001;
parameter [15:0] HANN_C391 = 16'b0011100111101001;
parameter [15:0] HANN_C392 = 16'b0011100100100000;
parameter [15:0] HANN_C393 = 16'b0011100001011000;
parameter [15:0] HANN_C394 = 16'b0011011110010000;
parameter [15:0] HANN_C395 = 16'b0011011011001001;
parameter [15:0] HANN_C396 = 16'b0011011000000001;
parameter [15:0] HANN_C397 = 16'b0011010100111011;
parameter [15:0] HANN_C398 = 16'b0011010001110100;
parameter [15:0] HANN_C399 = 16'b0011001110101110;
parameter [15:0] HANN_C400 = 16'b0011001011101001;
parameter [15:0] HANN_C401 = 16'b0011001000100100;
parameter [15:0] HANN_C402 = 16'b0011000101100000;
parameter [15:0] HANN_C403 = 16'b0011000010011100;
parameter [15:0] HANN_C404 = 16'b0010111111011001;
parameter [15:0] HANN_C405 = 16'b0010111100010110;
parameter [15:0] HANN_C406 = 16'b0010111001010100;
parameter [15:0] HANN_C407 = 16'b0010110110010011;
parameter [15:0] HANN_C408 = 16'b0010110011010010;
parameter [15:0] HANN_C409 = 16'b0010110000010010;
parameter [15:0] HANN_C410 = 16'b0010101101010011;
parameter [15:0] HANN_C411 = 16'b0010101010010101;
parameter [15:0] HANN_C412 = 16'b0010100111011000;
parameter [15:0] HANN_C413 = 16'b0010100100011011;
parameter [15:0] HANN_C414 = 16'b0010100001011111;
parameter [15:0] HANN_C415 = 16'b0010011110100101;
parameter [15:0] HANN_C416 = 16'b0010011011101011;
parameter [15:0] HANN_C417 = 16'b0010011000110010;
parameter [15:0] HANN_C418 = 16'b0010010101111010;
parameter [15:0] HANN_C419 = 16'b0010010011000011;
parameter [15:0] HANN_C420 = 16'b0010010000001101;
parameter [15:0] HANN_C421 = 16'b0010001101011001;
parameter [15:0] HANN_C422 = 16'b0010001010100101;
parameter [15:0] HANN_C423 = 16'b0010000111110011;
parameter [15:0] HANN_C424 = 16'b0010000101000001;
parameter [15:0] HANN_C425 = 16'b0010000010010001;
parameter [15:0] HANN_C426 = 16'b0001111111100010;
parameter [15:0] HANN_C427 = 16'b0001111100110101;
parameter [15:0] HANN_C428 = 16'b0001111010001000;
parameter [15:0] HANN_C429 = 16'b0001110111011101;
parameter [15:0] HANN_C430 = 16'b0001110100110100;
parameter [15:0] HANN_C431 = 16'b0001110010001011;
parameter [15:0] HANN_C432 = 16'b0001101111100100;
parameter [15:0] HANN_C433 = 16'b0001101100111111;
parameter [15:0] HANN_C434 = 16'b0001101010011010;
parameter [15:0] HANN_C435 = 16'b0001100111111000;
parameter [15:0] HANN_C436 = 16'b0001100101010110;
parameter [15:0] HANN_C437 = 16'b0001100010110111;
parameter [15:0] HANN_C438 = 16'b0001100000011000;
parameter [15:0] HANN_C439 = 16'b0001011101111100;
parameter [15:0] HANN_C440 = 16'b0001011011100000;
parameter [15:0] HANN_C441 = 16'b0001011001000111;
parameter [15:0] HANN_C442 = 16'b0001010110101111;
parameter [15:0] HANN_C443 = 16'b0001010100011001;
parameter [15:0] HANN_C444 = 16'b0001010010000100;
parameter [15:0] HANN_C445 = 16'b0001001111110001;
parameter [15:0] HANN_C446 = 16'b0001001101100000;
parameter [15:0] HANN_C447 = 16'b0001001011010000;
parameter [15:0] HANN_C448 = 16'b0001001001000010;
parameter [15:0] HANN_C449 = 16'b0001000110110110;
parameter [15:0] HANN_C450 = 16'b0001000100101100;
parameter [15:0] HANN_C451 = 16'b0001000010100100;
parameter [15:0] HANN_C452 = 16'b0001000000011101;
parameter [15:0] HANN_C453 = 16'b0000111110011000;
parameter [15:0] HANN_C454 = 16'b0000111100010101;
parameter [15:0] HANN_C455 = 16'b0000111010010100;
parameter [15:0] HANN_C456 = 16'b0000111000010101;
parameter [15:0] HANN_C457 = 16'b0000110110011000;
parameter [15:0] HANN_C458 = 16'b0000110100011101;
parameter [15:0] HANN_C459 = 16'b0000110010100100;
parameter [15:0] HANN_C460 = 16'b0000110000101101;
parameter [15:0] HANN_C461 = 16'b0000101110111000;
parameter [15:0] HANN_C462 = 16'b0000101101000100;
parameter [15:0] HANN_C463 = 16'b0000101011010011;
parameter [15:0] HANN_C464 = 16'b0000101001100100;
parameter [15:0] HANN_C465 = 16'b0000100111110111;
parameter [15:0] HANN_C466 = 16'b0000100110001100;
parameter [15:0] HANN_C467 = 16'b0000100100100011;
parameter [15:0] HANN_C468 = 16'b0000100010111101;
parameter [15:0] HANN_C469 = 16'b0000100001011000;
parameter [15:0] HANN_C470 = 16'b0000011111110110;
parameter [15:0] HANN_C471 = 16'b0000011110010110;
parameter [15:0] HANN_C472 = 16'b0000011100110111;
parameter [15:0] HANN_C473 = 16'b0000011011011100;
parameter [15:0] HANN_C474 = 16'b0000011010000010;
parameter [15:0] HANN_C475 = 16'b0000011000101011;
parameter [15:0] HANN_C476 = 16'b0000010111010101;
parameter [15:0] HANN_C477 = 16'b0000010110000011;
parameter [15:0] HANN_C478 = 16'b0000010100110010;
parameter [15:0] HANN_C479 = 16'b0000010011100011;
parameter [15:0] HANN_C480 = 16'b0000010010010111;
parameter [15:0] HANN_C481 = 16'b0000010001001110;
parameter [15:0] HANN_C482 = 16'b0000010000000110;
parameter [15:0] HANN_C483 = 16'b0000001111000001;
parameter [15:0] HANN_C484 = 16'b0000001101111110;
parameter [15:0] HANN_C485 = 16'b0000001100111110;
parameter [15:0] HANN_C486 = 16'b0000001100000000;
parameter [15:0] HANN_C487 = 16'b0000001011000100;
parameter [15:0] HANN_C488 = 16'b0000001010001010;
parameter [15:0] HANN_C489 = 16'b0000001001010011;
parameter [15:0] HANN_C490 = 16'b0000001000011111;
parameter [15:0] HANN_C491 = 16'b0000000111101100;
parameter [15:0] HANN_C492 = 16'b0000000110111101;
parameter [15:0] HANN_C493 = 16'b0000000110001111;
parameter [15:0] HANN_C494 = 16'b0000000101100100;
parameter [15:0] HANN_C495 = 16'b0000000100111100;
parameter [15:0] HANN_C496 = 16'b0000000100010101;
parameter [15:0] HANN_C497 = 16'b0000000011110010;
parameter [15:0] HANN_C498 = 16'b0000000011010000;
parameter [15:0] HANN_C499 = 16'b0000000010110010;
parameter [15:0] HANN_C500 = 16'b0000000010010101;
parameter [15:0] HANN_C501 = 16'b0000000001111011;
parameter [15:0] HANN_C502 = 16'b0000000001100100;
parameter [15:0] HANN_C503 = 16'b0000000001001111;
parameter [15:0] HANN_C504 = 16'b0000000000111100;
parameter [15:0] HANN_C505 = 16'b0000000000101100;
parameter [15:0] HANN_C506 = 16'b0000000000011110;
parameter [15:0] HANN_C507 = 16'b0000000000010011;
parameter [15:0] HANN_C508 = 16'b0000000000001011;
parameter [15:0] HANN_C509 = 16'b0000000000000100;
parameter [15:0] HANN_C510 = 16'b0000000000000001;
parameter [15:0] HANN_C511 = 16'b0000000000000000;